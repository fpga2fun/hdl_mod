sum = 81, val = 62 -20 39
sum = 39, val = -27 67 1 76 -97 -58 77
sum = 38, val = 60 -22
sum = 72, val =-120 29 123 102 -41 -21
sum = -53, val = -58 -85 -115 112 -101 -62