busif.cb.request <= 1;		//同步驱动
busif.cb.cmd <= cmd_buf;	//同步驱动