initital begin
 ascend = '{0,1,2,3};
 $display("%p",ascend); //'{0，1，2，3}
 ascend = '{4{8}};
 $display("%p",ascend); //'{8，8，8，8}
end