////////////////////////////////////////////////////////////////////
// Purpose: Top level testbench for Chap_6_Randomization/exercise11
// Author: Greg Tumbush
//
// REVISION HISTORY:
// $Log: top.sv,v $
// Revision 1.1  2011/05/29 19:09:54  tumbush.tumbush
// Check into cloud repository
//
// Revision 1.1  2011/05/10 20:10:55  Greg
// Initial check-in
//
/////////////////////////////////////////////////////////////////////
`default_nettype none
module top;

test test();
   
endmodule

