clocking cb @(posedge clk);
  output #10ns request;
  input #15ns grant;
endclocking
