bit [7:0] mask[] = '{
    8'b0000_0000,
    8'b0000_0001,
    8'b0000_0011,
    8'b0000_0111,
    8'b0000_1111,
    8'b0001_1111,
    8'b0011_1111,
    8'b0111_1111,
    8'b1111_1111
};
