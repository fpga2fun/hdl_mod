//////////////////////////////////////////////////////////////
// Purpose: Top level testbench for Chap_5_Basic_OOP/exercise6
// Author: Greg Tumbush
//
// REVISION HISTORY:
// $Log: top.sv,v $
// Revision 1.1  2011/05/29 19:03:49  tumbush.tumbush
// Check into cloud repository
//
// Revision 1.1  2011/05/09 13:31:18  Greg
// Initial check-in
//
/////////////////////////////////////////////////////////////
`default_nettype none
module top;

test test();
   
endmodule

