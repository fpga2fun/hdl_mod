##2 arbif.cb.request <= 0; // 等待两个时钟周期然后赋值
##3; // 非法 — 必须和赋值语句同时使用