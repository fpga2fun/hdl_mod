///////////////////////////////////////////////
// Purpose: DUT for Chap_2_Data_Types/exercise11
// Author: Greg Tumbush
//
// REVISION HISTORY:
// $Log: alu.v,v $
// Revision 1.1  2011/05/28 19:48:06  tumbush.tumbush
// Check into cloud repository
//
// Revision 1.1  2011/05/05 22:22:55  Greg
// Initial check-in
//
///////////////////////////////////////////////

`default_nettype none
  module alu(
    input wire [1:0] opcode
	     );
endmodule