sum = 1011, val = 83 249 197 187 152 95 40 8
sum = 1012, val = 213 252 213 44 196 20 20 54
sum = 370, val = 118 76 176
sum = 976, val = 233 187 44 157 201 81 73
sum = 412, val = 172 167 73