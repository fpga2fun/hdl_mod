lo = 20, med = 224, hi = 164
lo = 114, med = 39, hi = 189
lo = 186, med = 148, hi = 161
lo = 214, med = 223, hi = 201