a40: assert (arbif.cb.grant == 2'b01)
else $error("Grant not asserted");