task run();
  done = 0;
  while (!done) begin
    // 获取下一个事物
    // 进行变换
    // 发送事件
  end
endtask
