covergroup CovDst27;
  coverpoint tr.dst {
    ignore_bins hi = {6, 7};  // 忽略最后两个仓
  }
endgroup
