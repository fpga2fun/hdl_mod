typedef union { bit [31:0] b; int i; } num_u;
num_u un;
un.i = -1;// 把数值设为无符号整数