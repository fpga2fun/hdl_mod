int array2[0:7][0:3];  // 完整的声明
int array3[8][4];  // 紧凑的声明
array2[7][3] = 1;  // 设置最后一个元素
