class Xactor;
  task run();
    Print::error("NYI", "This Xactor is not yet implemented");
  endtask
endclass
