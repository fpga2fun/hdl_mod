sum = 79, val = 88 100 246 2 14 228 169
sum = 120, val = 74 75 141 86
sum = 39, val = 39
sum = 193, val = 31 156 172 33 57
sum = 173, val = 59 150 25 101 138 212