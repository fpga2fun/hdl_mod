typedef struct {bit [7:0] r, g, b;} pixel_s;
pixel_s my_pixel;
