class Driver;
  virtual X_if #(.BIT_WIDTH(BIT_WIDTH)) xi;
  //...
endclass
