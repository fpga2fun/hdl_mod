task automatic sticky(ref int array[50],
 input int a, b); // 明确指定方向