class Driver;
  vx_if xi;
  int   id;
  function new(input vx_if xi, input int id);
    this.xi = xi;
    this.id = id;
  endfunction
  //...
endclass : Driver
