import "DPI-C" function int addmul(
  input int a,
  b,
  output int sum
);
import "DPI-C" function void stop_model();
