import "DPI-C" pure function int factorial(input int i);
import "DPI-C" pure function real sin(input real in);
