covergroup CovDst25;
  coverpoint tr.dst {bins t1 = (0 => 1), (0 => 2), (0 => 3);}
endgroup
