////////////////////////////////////////////////////////////////////////////////
// Purpose: AHB slave for Chap_4_Connecting_the_Testbench_and_Design/exercise1
// Author: Greg Tumbush
//
// REVISION HISTORY:
// $Log: ahb_slave.sv,v $
// Revision 1.1  2011/05/28 20:22:55  tumbush.tumbush
// Check into cloud repository
//
// Revision 1.1  2011/05/08 22:13:59  Greg
// Initial check-in
//
////////////////////////////////////////////////////////////////////////////////
`default_nettype none
  module ahb_slave(ahb_if ahb_bus);
endmodule // ahb_slave
