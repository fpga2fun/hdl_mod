function void create(ref Transaction tr);
...
endfunction : create