logic [7:0] local_addr
local_addr = addr << 2; // 漏洞