task sticky(int a, b);