program automatic initialization; // 漏洞被修复
...
endprogram