program automatic test;
  import abc::*;
  Transaction tr;
  // 测试代码
endprogram
