class LogImp;
  rand bit d, e;
  constraint c {(d == 1) -> (e == 1);}
endclass
