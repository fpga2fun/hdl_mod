typedef union packed {
  uniType uni;
  nniType nni;
  bit [0:52][7:0] Mem;
} ATMCellType;
