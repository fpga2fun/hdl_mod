//////////////////////////////////////////////////////////////
// Purpose: Top level testbench for Chap_5_Basic_OOP/exercise7
// Author: Greg Tumbush
//
// REVISION HISTORY:
// $Log: top.sv,v $
// Revision 1.2  2011/07/21 23:32:15  tumbush.tumbush
// Replaced PrintBase with PrintUtilities. Converted with dos2unix.
//
// Revision 1.1  2011/05/09 13:35:23  Greg
// Initial check-in
//
/////////////////////////////////////////////////////////////
`default_nettype none
module top;

test test();
   
endmodule

