////////////////////////////////////////////////////////////////////
// Purpose: Top level testbench for Chap_6_Randomization/exercise5
// Author: Greg Tumbush
//
// REVISION HISTORY:
// $Log: top.sv,v $
// Revision 1.1  2011/05/29 19:09:59  tumbush.tumbush
// Check into cloud repository
//
// Revision 1.1  2011/05/10 18:55:32  Greg
// Initial check-in
//
/////////////////////////////////////////////////////////////////////
`default_nettype none
module top;

test test();
   
endmodule

