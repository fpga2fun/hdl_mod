C: in c_display
SV: In top.b1.sv_display
C: in c_display
SV: In top.sv_display