task mytask2 (output logic [31:0] x,
 input logic y);
...
endtask