typedef enum {
  FIRST  = 1,
  SECOND,
  THIRD
} ordinal_e;
ordinal_e position;
