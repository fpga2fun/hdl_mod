"test.sv", 7: top.t1.a1: started at 55ns failed at 55ns
offending '(arbif.cb.grant == 2'b1) '