module arb_with_mp (arb_if.DUT arbif);
 ...
endmodule