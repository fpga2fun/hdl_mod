Coverpoint Coverage report
CoverageGroup: CovDst2
 Coverpoint: tr.dst
Summary
 Coverage: 87.50
 Goal: 100
 Number of Expected auto-bins: 8
 Number of User Defined Bins: 0
 Number of Automatically Generated Bins: 7
 Number of User Defined Transitions: 0
 
 Automatically Generated Bins
 Bin # hits at least
 ================================
 auto[1] 7 1
 auto[2] 7 1
 auto[3] 1 1
 auto[4] 5 1
 auto[5] 4 1
 auto[6] 2 1
 auto[7] 6 1
 ================================