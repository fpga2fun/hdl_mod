Bin # hits at least
======================================
auto[0:3] 15 1
auto[4:7] 17 1
======================================