constraint c_fibonacci {
  (f == vals[0]) ||  // f==1
  (f == vals[1]) ||  // f==2
  (f == vals[2]) ||  // f==3
  (f == vals[3]) ||  // f==5
  (f == vals[4]);  // f==8
}
