module uses_a_port(inout bit not_connected);
 ...
endmodule