int d[] = '{9,1,8,3,4,4};
d.reverse();  // '{4,4,3,8,1,9}
d.sort();     // '{1,3,4,4,8,9}
d.rsort();    // '{9,8,4,4,3,1}
d.shuffle();  // '{9,4,3,8,1,4}
