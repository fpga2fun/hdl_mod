program automatic test (
    bus_ifc bus
);
  initial $display(bus.data);  // 使用接口信号
endprogram
