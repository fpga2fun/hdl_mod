Transaction src, dst;
initial begin
  src = new();  // 创建第一个对象
  dst = src.copy();  // 复制对象
end
