import "DPI-C" context task call_sv(bit [31:0] data);
