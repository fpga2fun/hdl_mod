typedef bit [63:0] bit64_t;
bit64_t assoc[bit64_t], idx = 1;
