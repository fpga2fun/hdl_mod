struct {bit [7:0] r, g, b;} pixel;
