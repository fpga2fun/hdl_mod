C: in c_display
SV: in sv_display