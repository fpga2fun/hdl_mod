case( graduation_year ) inside // 注意 “inside” 关键字
 [ 1950:1959 ]:$display ( "Do you like bobby sox? " );
 [ 1960:1969 ]:$display ( "Did you go to Woodstock? " );
 [ 1970:1979 ]:$display ( "Did you dance to disco? " );
endcase