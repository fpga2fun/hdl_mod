module atm_router(Rx_if.DUT Rx0, Rx1, Rx2, Rx3,
 Tx_if.DUT Tx0, Tx1, Tx2, Tx3,
 input logic clk, rst);
 ...
endmodule