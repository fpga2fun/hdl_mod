sum = 989, val = 787 202
sum = 1021, val = 564 76 132 235 0 8 6
sum = 872, val = 624 101 136 11
sum = 978, val = 890 88
sum = 905, val = 663 242