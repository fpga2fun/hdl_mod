// 文件 abc.svh
package abc;
  class Transaction;
    // 类主体
  endclass
endpackage
