typedef enum {
  INIT,
  DECODE = 2,
  IDLE
} fsmtype_e;
