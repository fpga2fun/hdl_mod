if ($isunknown(iport)==1)
$display("@%0t: 4-state value detected on iport %b",/
$time, iport);
