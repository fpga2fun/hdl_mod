Cumulative report for Transaction::CovDst30
Summary:
 Coverage: 78.91
 Goal: 100
Coverpoint Coverage Goal Weight
========================================================
kind 100.00 100 1
dst 100.00 100 1
========================================================
Cross Coverage Goal Weight
========================================================
Transaction::CovDst30 78.91 100 1
Cross Coverage report
CoverageGroup: Transaction::CovDst30
 Cross: Transaction::CovDst30
Summary
 Coverage: 36.72
 Goal: 100
 Coverpoints Crossed: kind dst
 Number of Expected Cross Bins: 128
 Number of User Defined Cross Bins: 0
 Number of Automatically Generated Cross Bins: 47
 Automatically Generated Cross Bins
 kind dst # hits at least
==================================================
auto[0] auto[0] 1 1
auto[0] auto[1] 2 1
auto[0] auto[2] 1 1
auto[0] auto[5] 1 1
...