tq = d.find_first with (item == 4);  // 本例的四个语句都是等价的
tq = d.find_first() with (item == 4);
tq = d.find_first(item) with (item == 4);
tq = d.find_first(x) with (x == 4);
