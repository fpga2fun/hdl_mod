mailbox #(Transaction) mbx_tr;  // 参数化信箱：建议的方式
mailbox mbx_untyped;  // 不专业：不建议
