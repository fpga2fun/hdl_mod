int f[6] = '{1, 6, 2, 6, 8, 6};  // 定宽数组
int d[] = '{2, 4, 6, 8, 10};  // 动态数组
int
    q[$] = {1, 3, 5, 7},  // 队列
    tq[$];  // 用来保存结果的临时队列
tq = q.min();  //{1}
tq = d.max();  //{10}
tq = f.unique();  //{1，6，2，8}
