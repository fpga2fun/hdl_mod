enum {
  RED,
  BLUE,
  GREEN
} color;
