a = $urandom_range(3, 10);  // 值的范围是 3-10
a = $urandom_range(10, 3);  // 值的范围是 3-10
b = $urandom_range(5);  // 值的范围是 0-5
