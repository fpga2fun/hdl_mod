M 100
W 12 34
W 99 8
R 12 34