int i;
real r;
i = int'(10.0 - 0.1);  // 转换是非强制的
r = real'(42);  // 转换是非强制的
