bit b;  // 双状态，单比特
bit [31:0] b32;  // 双状态，32 比特无符号整数
int unsigned ui;  // 双状态，32 比特无符号整数
int i;  // 双状态，32 比特有符号整数
byte b8;  // 双状态，8 比特有符号整数
shortint s;  // 双状态，16 比特有符号整数
longint l;  // 双状态，64 比特有符号整数
integer i4;  // 四状态，32 比特有符号整数
time t;  // 四状态，64 比特无符号整数
real r;  // 双状态，双精度浮点数
