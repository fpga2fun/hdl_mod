initial begin
  int h;
  bit [7:0] b, g[4], j[4] = '{8'ha, 8'hb, 8'hc, 8'hd};
  bit [7:0] q, r, s, t;
  h = {>>{j}};  //0a0b0c0d 把数组打包成整型
  h = {<<{j}};  //b030d050 位倒序
  h = {<<byte{j}};  //0d0c0b0a 字节倒序
  {>>{g}} = {<<byte{j}};  //0d，0c，0b，0a 拆分成数组
  b = {<<{8'b0011_0101}};  //1010_1100 位倒序
  b = {<<4{8'b0011_0101}};  //0101_0011 半字节倒序
  {>>{q, r, s, t}} = j;  // 把 j 分散到四个字节变量里
  h = {>>{t, s, r, q}};  // 把字节集中到 h 里
end
