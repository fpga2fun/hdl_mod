@0: 1: before trigger
@0: 2: before trigger
@0: 1: after trigger