#!/usr/local/bin/perl
print "Perl: Hello world!\n" ;
exit (3)