void'($fscanf(file, "%d", i));
