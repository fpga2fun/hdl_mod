////////////////////////////////////////////////////////////////////
// Purpose: Class definitions for Chap_6_Randomization/exercise4
// Author: Greg Tumbush
//
// REVISION HISTORY:
// $Log: top.sv,v $
// Revision 1.1  2011/05/29 19:09:57  tumbush.tumbush
// Check into cloud repository
//
// Revision 1.1  2011/05/10 18:19:35  Greg
// Initial check-in
//
/////////////////////////////////////////////////////////////////////
`default_nettype none
module top;

test test();
   
endmodule

