Transaction tr;  // 声明一个句柄
tr = new();  // 为一个 Transaction 对象分配空间
