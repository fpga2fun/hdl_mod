typedef enum {
  BAD_O  = 0,
  FIRST  = 1,
  SECOND,
  THIRD
} ordinal_e;
ordinal_e position;
