interface X_if (
    input logic clk
);
  // …
endinterface
typedef virtual X_if.TB vx_if;
