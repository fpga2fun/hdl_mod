////////////////////////////////////////////////////////////////////////////////////////
// Purpose: Testbench for Chap_7_Threads_and_Interprocess_Communication/homework2_solution
// Author: Greg Tumbush
//
// REVISION HISTORY:
// $Log: top.sv,v $
// Revision 1.1  2011/05/29 19:13:51  tumbush.tumbush
// Check into cloud repository
//
// Revision 1.1  2011/03/19 14:44:10  Greg
// Initial check in
//
/////////////////////////////////////////////////////////////////////////////////////////
`default_nettype none
module top;

test test();   

   
endmodule

