covergroup CovDst42;
  type_option.comment = "Section 3.2.14 Dst Port numbers";
  coverpoint tr.dst;
endgroup
