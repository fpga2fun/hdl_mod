C: c_display called from top.b1
C: Calling top.b1.sv_display
SV: In top.b1.sv_display
C: c_display called from top
C: Calling top.b1.sv_display
SV: In top.b1.sv_display