typedef bit [31:0] uint;  // 32 比特双状态无符号数
typedef int unsigned uint;  // 等效的定义
