covergroup CovDst29;
  coverpoint tr.dst {
    illegal_bins hi = {6, 7};  // 如果出现便报错
  }
endgroup
