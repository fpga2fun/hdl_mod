M 100