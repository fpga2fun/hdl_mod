covergroup CoverLength(ref bit [2:0] len);
  coverpoint len;
  option.per_instance = 1;
endgroup
