function bit transmit(input bit [31:0] data);
 // 发送处理
 ...
 return status; // 返回状态：0 = error
endfunction