`default_nettype none
module top;

test test();   

   
endmodule

