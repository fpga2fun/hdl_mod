covergroup CrossManual;
  ab: coverpoint {
    sam.a, sam.b
  } {
    bins a0b0 = {2'b00}; bins a1b0 = {2'b10}; wildcard bins b1 = {2'b?1};
  }
endgroup
