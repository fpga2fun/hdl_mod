covergroup CovDst12;
  coverpoint tr.dst {option.auto_bin_max = 2;}  // 分成 2 个仓
endgroup
