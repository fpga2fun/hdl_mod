virtual class svm_object;
  // 空类
endclass
