extern void sv_display();

void c_display() {
 io_printf("C: in c_display\n");
 sv_display();
}