covergroup CovDst45;
  coverpoint tr.dst;
  option.goal = 90;  // 只需要部分覆盖即可满足
endgroup
