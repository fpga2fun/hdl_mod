////////////////////////////////////////////////////////////////////
// Purpose: Top level testbench for Chap_6_Randomization/exercise1_3
// Author: Greg Tumbush
//
// REVISION HISTORY:
// $Log: top.sv,v $
// Revision 1.1  2011/05/29 19:09:55  tumbush.tumbush
// Check into cloud repository
//
// Revision 1.1  2011/05/10 16:20:24  Greg
// Initial check-in
//
/////////////////////////////////////////////////////////////////////
`default_nettype none
module top;

test test();
   
endmodule

