typedef class Statistics; // 定义低级别类

class Transaction;
 Statistics stats; // 使用 Statistics 类
 ...
endclass

class Statistics; // 定义 Statistics 类
 ...
endclass