constraint c_range {
  !(c inside {[lo : hi]});  // c < lo 或 c > hi
}
