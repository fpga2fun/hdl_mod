//////////////////////////////////////////////////////////////////////////
// Purpose: SystemVerilog module for Chap_12_Interfacing_with_C/exercise7
// Author: Chris Spear
//
// REVISION HISTORY:
// $Log: top.sv,v $
// Revision 1.2  2011/09/27 17:21:37  tumbush.tumbush
// Added header information
//
//
//////////////////////////////////////////////////////////////////////////
module top;

   test test();
   
endmodule // top
