task T3;
    input a, b;
    logic a, b;
    output [15:0] u, v;
    bit [15:0] u, v;
    ...
endtask
