int lo_hi[0:15];  // 16 个整数 [0]..[15]
int c_style[16];  // 16 个整数 [0]..[15]
