/////////////////////////////////////////////////////////////////
// Purpose: Top level testbench for Chap_6_Randomization/exercise9
// Author: Greg Tumbush
//
// REVISION HISTORY:
// $Log: top.sv,v $
// Revision 1.1  2011/05/29 19:10:03  tumbush.tumbush
// Check into cloud repository
//
// Revision 1.1  2011/05/10 19:56:06  Greg
// Initial check-in
//
/////////////////////////////////////////////////////////////////

`default_nettype none
module top;

test test();
   
endmodule

