//////////////////////////////////////////////////////////////
// Purpose: Top level testbench for Chap_5_Basic_OOP/exercise4
// Author: Greg Tumbush
//
// REVISION HISTORY:
// $Log: top.sv,v $
// Revision 1.1  2011/05/29 19:03:46  tumbush.tumbush
// Check into cloud repository
//
// Revision 1.1  2011/05/09 13:23:06  Greg
// Initial check-in
//
/////////////////////////////////////////////////////////////
`default_nettype none
module top;

test test();
   
endmodule

