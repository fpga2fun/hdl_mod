package ABC;
  parameter int abc_data_width = 32;
  typedef logic [abc_data_width-1:0] abc_data_t;
  parameter time timeout = 100ns;
  string message = "ABC done";
endpackage  //ABC
