//////////////////////////////////////////////////////////////
// Purpose: Package for Chap_5_Basic_OOP/exercise8
// Author: Greg Tumbush
//
// REVISION HISTORY:
// $Log: my_package.sv,v $
// Revision 1.1  2011/05/29 19:03:51  tumbush.tumbush
// Check into cloud repository
//
// Revision 1.1  2011/05/09 13:40:12  Greg
// Initial check-in
//
/////////////////////////////////////////////////////////////
package automatic my_package;
   
class Transaction;	
   logic [7:0] addr;
endclass // Transaction

  endpackage
