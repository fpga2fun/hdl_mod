task mytask1;
 output [31:0] x;
 reg [31:0] x;
 input y;
 ...
endtask