virtual class svm_object_wrapper;
  pure virtual function string get_type_name();
  pure virtual function svm_object create_object(string name);
endclass
