/////////////////////////////////////////////////////////////////////////////////
// Purpose: Top for Chap_7_Threads_and_Interprocess_Communication/exercise4_5
// Author: Chris Spear
//
// REVISION HISTORY:
// $Log: top.sv,v $
// Revision 1.1  2011/05/29 19:13:45  tumbush.tumbush
// Check into cloud repository
//
// Revision 1.1  2011/05/10 23:17:52  Greg
// Initial check-in
//
/////////////////////////////////////////////////////////////////////////////////
`default_nettype none
module top;

test test();
   
endmodule

