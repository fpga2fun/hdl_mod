Summary
 Coverage: 90.91
 Number of Coverpoints Crossed: 2
 Coverpoints Crossed: kind dst
 Number of Expected Cross Bins: 88
 Number of Automatically Generated Cross Bins: 80
 Automatically Generated Cross Bins
 dst kind # hits at least
 ======================================================
 dst_0 hi_8 3 1
 dst_0 hi_a 1 1
 dst_0 hi_b 4 1
 dst_0 hi_c 4 1
 dst_0 hi_d 4 1
 dst_0 hi_e 1 1
 dst_0 lo 7 1
 dst_0 zero 1 1
 dst_1 hi_8 3 1