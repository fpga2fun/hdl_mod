//////////////////////////////////////////////////////////////////////
// Purpose: Top level module for Chap_12_Interfacing_with_C/exercise4_slide
// Author: Greg Tumbush
//
// REVISION HISTORY:
// $Log: top.sv,v $
// Revision 1.1  2011/09/27 19:43:57  tumbush.tumbush
// Initial check-in
//
//
//////////////////////////////////////////////////////////////////////
module top;

   test test();
   
endmodule // top
