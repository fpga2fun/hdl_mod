driver drv;
drv = driver::type_id::create("drv", this);
