Bin # hits at least
============================
len_00 13 1
len_01 36 1
len_02 51 1
len_03 60 1
len_04 72 1
len_05 88 1
len_06 127 1
len_07 122 1
len_08 133 1
len_09 138 1
len_0a 115 1
len_0b 128 1
len_0c 125 1
len_0d 111 1
len_0e 115 1
len_0f 134 1
len_10 107 1
len_11 102 1
len_12 70 1
len_13 65 1
len_14 39 1
len_15 30 1
len_16 19 1
len_17 0 1
============================