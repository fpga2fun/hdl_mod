sum = 245, val = 1348956995 3748256598 985546882 2507174362
sum = 600, val = 2072193829 315191491 484497976 3050698208
 2300168220 3988671456 3998079060 970369544
sum = 17, val = 1924767007 3550820640 4149215303 3260098955
sum = 440, val = 3192781444 624830067 1300652226 4072252356
 3694386235
sum = 864, val = 3561488468 733479692