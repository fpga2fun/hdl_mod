> simv + script = ”perl hellp.pl”