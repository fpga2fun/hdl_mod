program automatic test #(
    NUM_XI = 2
);
  vx_if vxi[NUM_XI];  // 虚拟接口数组
  Driver driver[];
  //...
endprogram
