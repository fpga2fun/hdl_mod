byte b[$] = {2, 3, 4, 5};
int w;
w = b.sum();  // 14 = 2 + 3 + 4 + 5
w = b.product();  //120 = 2 * 3 * 4 * 5
w = b.and();  //0000_0000 = 2 & 3 & 4 & 5
