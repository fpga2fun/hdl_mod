"test.sv", 7: top.t1.a40: started at 55ns failed at 55ns
Offending '(arbif.cb.grant == 2'b01)'
Error: "test.sv", 7: top.t1.a40: at time 55 ns
Grant not asserted