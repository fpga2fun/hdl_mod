Transaction t; // 声明一个 Transaction 句柄
t = new(); // 创建一个 Transaction 对象
t.addr = 32'h42; // 设置变量的值
t.display(); // 调用一个子程序