task automatic sticky(ref int array[50],
 int a, b); // 这些参数的方向是什么？