initial begin
 const byte colon = ":";
 ...
end