covergroup CovDst44;
 kind: coverpoint tr.kind;
 dst: coverpoint tr.dst
 cross kind, dst;
 option.cross_num_print_missing = 1_000;
endgroup