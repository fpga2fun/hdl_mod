import "DPI-C" function chandle counter7_new();
import "DPI-C" function void counter7(
  input chandle inst,
  output logic [6:0] out,
  input logic [6:0] in,
  input logic reset,
  load
);
