////////////////////////////////////////////////////////////////////////////////////////////
// Purpose: Top level testbench for Chap_8_Advanced_OOP_and_Testbench_Guidelines/exercise5
// Author: Greg Tumbush
//
// REVISION HISTORY:
// $Log: top.sv,v $
// Revision 1.1  2011/05/29 19:16:06  tumbush.tumbush
// Check into cloud repository
//
// Revision 1.1  2011/05/11 22:40:05  Greg
// Initial check-in
//
////////////////////////////////////////////////////////////////////////////////////////////
`default_nettype none
module top;

test test();   

   
endmodule

