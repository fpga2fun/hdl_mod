Bin # hits at least
==================================
auto_DECODE 11 1
auto_IDLE 11 1
auto_INIT 10 1
==================================