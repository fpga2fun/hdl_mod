count[1]= 3980 ***************************************
count[2]= 3924 **************************************
count[3]= 3922 **************************************
count[5]= 4175 *****************************************
count[8]= 3999 ***************************************