module test_with_mp (arb_if.TEST arbif);
 ...
endmodule