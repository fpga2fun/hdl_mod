bit [7:0] b_unpack[3];  // 非合并数组
