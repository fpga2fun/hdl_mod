task multiple_lines;
  $display("First line");
  $display("Second line");
endtask : multiple_lines
