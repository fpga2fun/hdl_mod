////////////////////////////////////////////////////////////////////
// Purpose: Top level testbench for Chap_6_Randomization/exercise10
// Author: Greg Tumbush
//
// REVISION HISTORY:
// $Log: top.sv,v $
// Revision 1.1  2011/05/29 19:09:53  tumbush.tumbush
// Check into cloud repository
//
// Revision 1.1  2011/05/10 20:04:07  Greg
// Initial check-in
//
/////////////////////////////////////////////////////////////////////
`default_nettype none
module top;

test test();
   
endmodule

