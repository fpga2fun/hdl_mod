int
    j = 1,
    q2[$] = {3, 4},  // 队列的常量不需要使用 “'”
    q[$] = {0, 2, 5};  // {0,2,5}

initial begin  // 结果
  q = {q[0], j, q[1:$]};  // {0,1,2,5}     在 2 之前插入 1
  q = {q[0:2], q2, q[3:$]};  // {0,1,2,3,4,5}   在 q 中插入一个队列
  q = {q[0], q[2:$]};  // {0,2,3,4,5}   删除第 1 个元素

  // 下面的操作执行速度很快
  q = {6, q};  // {6,0,2,3,4,5} 在队列前面插入

  j = q[$];  //j = 5   从队列末尾取出数据
  q = q[0:$-1];  // {6,0,2,3,4}   效果和上一行相同

  q = {q, 8};  // {6,0,2,3,4,8} 在队列末尾插入

  j = q[0];  //j = 6   从队列前面取出数据
  q = q[1:$];  // {0,2,3,4,8}   效果和上一行相同

  q = {};  // {}   清空队列
end
